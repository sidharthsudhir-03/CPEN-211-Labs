module lab7_top(KEY,SW,LEDR,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5); 

	input[3:0]KEY; 
	input[9:0]SW; 
	output[9:0]LEDR; 
	output[6:0]HEX0,HEX1,HEX2,HEX3,HEX4,HEX5;
	
endmodule



