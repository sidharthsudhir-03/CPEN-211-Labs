module tb_lab3();

endmodule: tb_lab3
