module datapath_tb();

endmodule:datapath_tb