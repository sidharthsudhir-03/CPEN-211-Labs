module datapath();

endmodule:datapath