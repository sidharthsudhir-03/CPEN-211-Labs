module shifter_tb();

endmodule:shifter_tb