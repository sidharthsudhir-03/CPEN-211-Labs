module tb_lab3_gate();

endmodule: tb_lab3_gate
