module regfile_tb();

endmodule: regfile_tb