module ALU_tb();

endmodule: ALU_tb